--***************************************
--* TITLE: PNGenerator (receiver)	*
--* TYPE: Component 			*
--* AUTHOR: Dylan Van Assche 		*
--* DATE: 29/11/2017 			*
--***************************************
--* DESCRIPTION *
--***************
--1)Purpose:
-- Generating a PN code to match with the sender
--2)Principle:
-- Lineair feedback register to generate a PN code (31 bits) 
-- and which is restarted as soon a a PN code is found by the Matched Filter.
-- When the whole PN code is generated by the PN Generator a full_seq is 
-- triggered which is the bitsample signal (bit is ready for sampling).
--3)Inputs:
-- seq_det, rst, clk, clk_en
--4)Outputs:
-- full_seq, pn_1, pn_2, pn_3
--**********************
--* LIBRARIES & ENTITY *
--**********************
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
ENTITY pngenerator IS
PORT
(
	clk        : IN std_logic;
	clk_en     : IN std_logic;
	rst        : IN std_logic;
	seq_det    : IN std_logic;
	chipsample : IN std_logic;
	bitsample  : OUT std_logic;
	pn_1       : OUT std_logic;
	pn_2       : OUT std_logic;
	pn_3       : OUT std_logic
);
END;
--*********************************************
--* ARCHITECTURE, SIGNALS, TYPES & COMPONENTS *
--*********************************************
ARCHITECTURE behavior OF pngenerator IS
	SIGNAL shdata1          : std_logic_vector(4 DOWNTO 0) := "00010";
	SIGNAL shdata1_next     : std_logic_vector(4 DOWNTO 0) := (OTHERS => '0');
	SIGNAL shdata2          : std_logic_vector(4 DOWNTO 0) := "00111";
	SIGNAL shdata2_next     : std_logic_vector(4 DOWNTO 0) := (OTHERS => '0');
	SIGNAL full_seq_next    : std_logic;
	SIGNAL full_seq         : std_logic := '0';
	SIGNAL linear_feedback1 : std_logic := '0';
	SIGNAL linear_feedback2 : std_logic := '0';
BEGIN
-- calculate linear feedback for both PN counters (LFSR)
linear_feedback1 <= (shdata1(0) XOR shdata1(3));
linear_feedback2 <= ((shdata2(0) XOR shdata2(1)) XOR shdata2(3)) XOR shdata2(4);
-- connect signals to outputs
pn_1 <= shdata1(0);
pn_2 <= shdata2(0);
pn_3 <= shdata1(0) XOR shdata2(0);
bitsample <= full_seq;
-- 2-Process: synchronous part
pn_sync : PROCESS (clk)
BEGIN
	IF (rising_edge(clk) AND clk_en = '1' AND chipsample = '1') THEN
		IF (rst = '1') THEN -- rst line high, go to initial state
			shdata1 <= "00010"; -- constants aren't working here, signals become undefined
			shdata2 <= "00111";
			full_seq <= '0';
		ELSE -- normal operation
			full_seq <= full_seq_next;
			shdata1 <= shdata1_next;
			shdata2 <= shdata2_next;
		END IF;
	END IF;
END PROCESS pn_sync;
-- 2-Process: combinatoric part
pn_comb : PROCESS (shdata1, shdata2, linear_feedback1, linear_feedback2, seq_det, full_seq)
BEGIN
	IF (seq_det = '1') THEN
		shdata1_next <= "00010";
		shdata2_next <= "00111";
	ELSE
		shdata1_next <= linear_feedback1 & shdata1(4 DOWNTO 1);
		shdata2_next <= linear_feedback2 & shdata2(4 DOWNTO 1);
		IF (shdata1 = "00010") THEN -- next value is the "00001" value, prepare this already
			full_seq_next <= '1';
		ELSE
			full_seq_next <= '0';
		END IF;	
	END IF;
END PROCESS pn_comb;
END behavior;

